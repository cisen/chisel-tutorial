module VecShiftRegisterParam(
  input        clock,
  input        reset,
  input  [3:0] io_in,
  output [3:0] io_out
);
  assign io_out = 4'h0; // @[VecShiftRegisterParam.scala 20:10]
endmodule
