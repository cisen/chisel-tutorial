module VecShiftRegisterSimple(
  input        clock,
  input        reset,
  input  [7:0] io_in,
  output [7:0] io_out
);
  assign io_out = 8'h0; // @[VecShiftRegisterSimple.scala 22:10]
endmodule
