module Adder(
  input   clock,
  input   reset,
  input   io_in0,
  input   io_in1,
  output  io_out
);
  assign io_out = 1'h0; // @[Adder.scala 19:10]
endmodule
